`ifndef __DEFINES_SVH
`define __DEFINES_SVH

// ALU operands
`define     ALU_MOV     5'b00000
`define     ALU_ADD     5'b00001
`define     ALU_SUB     5'b00010
`define     ALU_AND     5'b00011
`define     ALU_OR      5'b00100
`define     ALU_NOT     5'b00101
`define     ALU_DEC     5'b00110
`define     ALU_INC     5'b00111
`define     ALU_MUL     5'b01000
`define     ALU_MOVU    5'b10000
`define     ALU_MOVL    5'b10100

`endif // __DEFINES_SVH