module RISC16(
);
    
endmodule // RISC16